/*
*
*	Creator : Ahmad Adel <github.com/ahmadadel8>
*						Dina  Elsokary <github.com/dinaelsokary>
*
* Contributer: Ahmad Hegazy <github.com/ahegazy> <ahegazipro@gmail.com>
*	Date: September 2018
* 
* Description: AddRoundKey step in AES encryption/Decryption.
* Language: Verilog
*
*/

module AddRoundKey
	#(parameter word_size =8 ,array_size =16)(
	input wire [word_size*array_size-1:0] key ,
	input wire [word_size*array_size-1:0] state,
	input  clk,enable, rst, load,
	output reg  [word_size*array_size-1:0]state_out,
	output reg done);
integer i,j,k,add;

task Mod;
	input  [14:0]x;
	output [7:0] y;

	reg    [8:0] con;
	reg    [14:0] z;
	integer i;
	 
	begin
		con = 9'd283;
		z = x;
		for (i=14; i>=8; i =i-1)
		 if (z > 8'd255)
			 begin
				if(z[i] == 1)
					z[i -: 9] = z[i -: 9] ^ con[8:0];
					//$display("z = %b",z[14:0]);
					end
		 else begin
			y =z;
			end
			y = z;
	end

endtask


always@(posedge clk)
 begin
 if (rst) begin
 state_out=128'd0;
 done <= 0;
 end 
 else if (enable) begin 
	for ( i=0; i<=15; i=i+1)
		Mod(key[i*word_size  +:  word_size] ^ state[i*word_size  +:  word_size],state_out[i*word_size  +:  word_size]);
////////////////////////////////////////////////
	done = 1;
end 
			else done <= 0;

end
endmodule

