class aes_configuration extends uvm_object;
	`uvm_object_utils(aes_configuration)

	function new(string name = "");
		super.new(name);
	endfunction: new
endclass: aes_configuration
